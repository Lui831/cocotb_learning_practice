-- simple_state_machine_pkg.vhd

library ieee;
use ieee.std_logic_1164.ALL;

-- Package initialziation
package simple_state_machine_pkg is
    
-- States of the state machine
type t_states is (RESET, IDLE, STATE1, STATE2, STATE3);



end simple_state_machine_pkg;

-- Package body
package body simple_state_machine_pkg is

end simple_state_machine_pkg;